netcdf bathymetry {
dimensions:
    x = 5;
    y = 5;

variables:
    double x(x);
        x:long_name = "X Coordinate";
        x:units = "meters";

    double y(y);
        y:long_name = "Y Coordinate";
        y:units = "meters";

    double z(y, x);
        z:long_name = "Bathymetry";
        z:units = "meters";

data:
    x = 0, 1, 2, 3, 4 ;
    y = 0, 1, 2, 3, 4 ;
    z =
        -20, -20, -20, -20, -20,      //Bathymetrievalues for y = 0
        -20, -30, -30, -30, -20,
        -20, -30, -40, -30, -20,
        -20, -30, -30, -30, -20,
        -20, -20, -20, -20, -20;      //Batymetrievalues for y = 4
}