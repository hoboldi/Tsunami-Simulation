netcdf displacment {
dimensions:
    x = 5;
    y = 5;

variables:
    double x(x);
        x:long_name = "X Coordinate";
        x:units = "meters";

    double y(y);
        y:long_name = "Y Coordinate";
        y:units = "meters";

    double z(y, x);
        z:long_name = "Displacement";
        z:units = "meters";

// global attributes:
                :Conventions = "COARDS" ;
data:
    x = 0, 1, 2, 3, 4 ;
    y = 0, 1, 2, 3, 4 ;
    z =
        0,0,0,0,0,
        -10,-10,-10,-10,-10,
        -20,-20,-20,-20,-20,
        -10, -10, -10, -10, -10,
        0,0,0,0,0 ;

}